package shared_pkg;

	int Error_count, Correct_count;
	bit test_finished;

endpackage